-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II"
-- VERSION		"Version 9.0 Build 132 02/25/2009 SJ Full Version"
-- CREATED ON		"Tue Jun 13 15:49:57 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY logicProcess IS 
	PORT
	(
		B0 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		B2 :  IN  STD_LOGIC;
		B3 :  IN  STD_LOGIC;
		B4 :  IN  STD_LOGIC;
		q1 :  IN  STD_LOGIC;
		q2 :  IN  STD_LOGIC;
		q3 :  IN  STD_LOGIC;
		q4 :  IN  STD_LOGIC;
		q5 :  IN  STD_LOGIC;
		q6 :  IN  STD_LOGIC;
		q7 :  IN  STD_LOGIC;
		q8 :  IN  STD_LOGIC;
		q9 :  IN  STD_LOGIC;
		q10 :  IN  STD_LOGIC;
		x1 :  OUT  STD_LOGIC;
		x2 :  OUT  STD_LOGIC;
		x3 :  OUT  STD_LOGIC;
		x4 :  OUT  STD_LOGIC;
		x5 :  OUT  STD_LOGIC;
		x6 :  OUT  STD_LOGIC;
		x7 :  OUT  STD_LOGIC;
		x8 :  OUT  STD_LOGIC;
		x9 :  OUT  STD_LOGIC;
		x10 :  OUT  STD_LOGIC;
		x11 :  OUT  STD_LOGIC;
		x12 :  OUT  STD_LOGIC;
		x13 :  OUT  STD_LOGIC;
		x14 :  OUT  STD_LOGIC;
		x15 :  OUT  STD_LOGIC;
		x16 :  OUT  STD_LOGIC;
		x17 :  OUT  STD_LOGIC;
		x18 :  OUT  STD_LOGIC
	);
END logicProcess;

ARCHITECTURE bdf_type OF logicProcess IS 

ATTRIBUTE black_box : BOOLEAN;
nATTRIBUTE noopt : BOOLEAN;

COMPONENT or5_0
	PORT(IN1 : IN STD_LOGIC;
		 IN3 : IN STD_LOGIC;
		 IN2 : IN STD_LOGIC;
		 IN5 : IN STD_LOGIC;
		 IN4 : IN STD_LOGIC;
		 OUT : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF or5_0: COMPONENT IS true;
ATTRIBUTE noopt OF or5_0: COMPONENT IS true;

COMPONENT logicpr2
	PORT(B0 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 B3 : IN STD_LOGIC;
		 B4 : IN STD_LOGIC;
		 L0 : OUT STD_LOGIC;
		 L1 : OUT STD_LOGIC;
		 L2 : OUT STD_LOGIC;
		 L3 : OUT STD_LOGIC;
		 L4 : OUT STD_LOGIC;
		 L5 : OUT STD_LOGIC;
		 L6 : OUT STD_LOGIC;
		 L7 : OUT STD_LOGIC;
		 L8 : OUT STD_LOGIC;
		 L9 : OUT STD_LOGIC;
		 L10 : OUT STD_LOGIC;
		 L11 : OUT STD_LOGIC;
		 L12 : OUT STD_LOGIC;
		 L13 : OUT STD_LOGIC;
		 L14 : OUT STD_LOGIC;
		 L15 : OUT STD_LOGIC;
		 L16 : OUT STD_LOGIC;
		 L17 : OUT STD_LOGIC;
		 L18 : OUT STD_LOGIC;
		 L19 : OUT STD_LOGIC;
		 L20 : OUT STD_LOGIC;
		 L21 : OUT STD_LOGIC;
		 L22 : OUT STD_LOGIC;
		 L23 : OUT STD_LOGIC;
		 L24 : OUT STD_LOGIC;
		 L25 : OUT STD_LOGIC;
		 L26 : OUT STD_LOGIC;
		 L27 : OUT STD_LOGIC;
		 L28 : OUT STD_LOGIC;
		 L29 : OUT STD_LOGIC;
		 L30 : OUT STD_LOGIC;
		 L31 : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;


BEGIN 
x3 <= SYNTHESIZED_WIRE_10;
x6 <= SYNTHESIZED_WIRE_17;
x11 <= SYNTHESIZED_WIRE_19;
x12 <= SYNTHESIZED_WIRE_20;
x13 <= SYNTHESIZED_WIRE_22;
x14 <= SYNTHESIZED_WIRE_21;
x17 <= SYNTHESIZED_WIRE_24;



b2v_inst : logicpr2
PORT MAP(B0 => B0,
		 B1 => B1,
		 B2 => B2,
		 B3 => B3,
		 B4 => B4,
		 L0 => SYNTHESIZED_WIRE_3,
		 L3 => SYNTHESIZED_WIRE_49,
		 L8 => x8,
		 L11 => SYNTHESIZED_WIRE_55,
		 L14 => SYNTHESIZED_WIRE_57,
		 L17 => SYNTHESIZED_WIRE_56,
		 L19 => SYNTHESIZED_WIRE_52,
		 L22 => SYNTHESIZED_WIRE_11,
		 L27 => SYNTHESIZED_WIRE_53);


b2v_inst1 : or5_0
PORT MAP(IN1 => SYNTHESIZED_WIRE_0,
		 IN3 => SYNTHESIZED_WIRE_1,
		 IN2 => SYNTHESIZED_WIRE_2,
		 IN5 => SYNTHESIZED_WIRE_3,
		 IN4 => SYNTHESIZED_WIRE_4,
		 OUT => x1);


SYNTHESIZED_WIRE_10 <= SYNTHESIZED_WIRE_49 OR SYNTHESIZED_WIRE_50 OR SYNTHESIZED_WIRE_7 OR SYNTHESIZED_WIRE_51;


x4 <= SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10;


SYNTHESIZED_WIRE_9 <= q9 AND SYNTHESIZED_WIRE_11;


SYNTHESIZED_WIRE_54 <= q3 AND SYNTHESIZED_WIRE_52;


SYNTHESIZED_WIRE_14 <= q9 AND SYNTHESIZED_WIRE_53;


x5 <= SYNTHESIZED_WIRE_14 OR SYNTHESIZED_WIRE_54;


SYNTHESIZED_WIRE_17 <= q1 AND SYNTHESIZED_WIRE_55;


SYNTHESIZED_WIRE_34 <= SYNTHESIZED_WIRE_17 OR SYNTHESIZED_WIRE_54 OR SYNTHESIZED_WIRE_19 OR SYNTHESIZED_WIRE_20 OR SYNTHESIZED_WIRE_21 OR SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_23 OR SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_55 AND q2;


SYNTHESIZED_WIRE_20 <= q4 AND SYNTHESIZED_WIRE_52;


SYNTHESIZED_WIRE_4 <= q3 AND SYNTHESIZED_WIRE_55;


SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_55 AND q5;


SYNTHESIZED_WIRE_21 <= SYNTHESIZED_WIRE_55 AND q6;


SYNTHESIZED_WIRE_23 <= SYNTHESIZED_WIRE_55 AND q7;


SYNTHESIZED_WIRE_24 <= SYNTHESIZED_WIRE_56 AND q8;


SYNTHESIZED_WIRE_33 <= q9 AND SYNTHESIZED_WIRE_53;


x7 <= SYNTHESIZED_WIRE_33 OR SYNTHESIZED_WIRE_34;


x9 <= SYNTHESIZED_WIRE_56 AND q10;


x10 <= SYNTHESIZED_WIRE_51 OR SYNTHESIZED_WIRE_50 OR SYNTHESIZED_WIRE_49;


x15 <= SYNTHESIZED_WIRE_55 AND q8;


x16 <= SYNTHESIZED_WIRE_57 AND q8;


SYNTHESIZED_WIRE_1 <= q4 AND SYNTHESIZED_WIRE_55;


x18 <= SYNTHESIZED_WIRE_55 AND q10;


SYNTHESIZED_WIRE_2 <= q9 AND SYNTHESIZED_WIRE_55;


SYNTHESIZED_WIRE_0 <= q10 AND SYNTHESIZED_WIRE_57;


x2 <= q9 AND SYNTHESIZED_WIRE_52;


SYNTHESIZED_WIRE_51 <= q3 AND SYNTHESIZED_WIRE_57;


SYNTHESIZED_WIRE_50 <= q4 AND SYNTHESIZED_WIRE_57;


SYNTHESIZED_WIRE_7 <= q9 AND SYNTHESIZED_WIRE_57;


END bdf_type;